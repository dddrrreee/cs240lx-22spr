module mux
    (
        input logic a, b,
        input logic sel,
        output logic out
    );
    // TODO
endmodule
