module adder
    (
        input logic [31:0] a, b,
        output logic [31:0] sum
    );
    // TODO
endmodule

module half_adder
    (
        input logic a, b,
        output logic c, s
    );
    // TODO
endmodule

module full_adder
    (
        input logic a, b, cin,
        output logic cout, s
    );
    // TODO
endmodule
